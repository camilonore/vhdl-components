library verilog;
use verilog.vl_types.all;
entity divisor_2_vlg_vec_tst is
end divisor_2_vlg_vec_tst;
