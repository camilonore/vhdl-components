library verilog;
use verilog.vl_types.all;
entity multiplicador_8_bits_vlg_vec_tst is
end multiplicador_8_bits_vlg_vec_tst;
