library verilog;
use verilog.vl_types.all;
entity multiplicador_4bits_vlg_vec_tst is
end multiplicador_4bits_vlg_vec_tst;
