library verilog;
use verilog.vl_types.all;
entity divisor_2_25_vlg_check_tst is
    port(
        oClk            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end divisor_2_25_vlg_check_tst;
