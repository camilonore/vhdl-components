library verilog;
use verilog.vl_types.all;
entity divisor_2 is
    port(
        Clk             : in     vl_logic;
        oClk            : out    vl_logic
    );
end divisor_2;
