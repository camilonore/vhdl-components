library verilog;
use verilog.vl_types.all;
entity restador_6bits_vlg_vec_tst is
end restador_6bits_vlg_vec_tst;
