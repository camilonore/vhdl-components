library verilog;
use verilog.vl_types.all;
entity bin_2_bcd_vlg_vec_tst is
end bin_2_bcd_vlg_vec_tst;
