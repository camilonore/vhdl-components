library ieee;
use ieee.std_logic_1164.all;

entity t_flipflop is
	port(
		T, R, P, Clk : in  std_logic := '0';
		       Q, nQ : out std_logic
	);
end t_flipflop;

architecture Behavioral of t_flipflop is
	
	signal tmp : std_logic := '0';
	
begin

	process(T, R, P, Clk) 
	
	begin
		if P = '1' then
			tmp <= '1';
		elsif R = '1' then
			tmp <= '0';
		elsif falling_edge(Clk) and T = '1' then 			
			tmp <= not(tmp);	
		elsif falling_edge(Clk) and T = '0' then 				
			tmp <= tmp;
		end if;	
	end process;
	
	Q  <= tmp;
	nQ <= not(tmp);
	
end Behavioral;
