library verilog;
use verilog.vl_types.all;
entity restador_4bits_vlg_vec_tst is
end restador_4bits_vlg_vec_tst;
