library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity bin_bcd is
	port ( 
	 Bin : in   std_logic_vector (7 downto 0);
	 Cen : out  std_logic_vector (3 downto 0);
	 Dec : out  std_logic_vector (3 downto 0);
	 Uni : out  std_logic_vector (3 downto 0)
	);
end bin_bcd;

architecture Behavioral of bin_bcd is

begin

    process(Bin)
        variable x: std_logic_vector (11 downto 0):= "000000000000";
    begin
	 
			
			if Bin = "00000000" then
			  x := "000000000000";
			elsif Bin = "00000001" then
			  x := "000000000001";
			elsif Bin = "00000010" then
			  x := "000000000010";
			elsif Bin = "00000011" then
			  x := "000000000011";
			elsif Bin = "00000100" then
			  x := "000000000100";
			elsif Bin = "00000101" then
			  x := "000000000101";
			elsif Bin = "00000110" then
			  x := "000000000110";
			elsif Bin = "00000111" then
			  x := "000000000111";
			elsif Bin = "00001000" then
			  x := "000000001000";
			elsif Bin = "00001001" then
			  x := "000000001001";
			elsif Bin = "00001010" then
			  x := "000000010000";
			elsif Bin = "00001011" then
			  x := "000000010001";
			elsif Bin = "00001100" then
			  x := "000000010010";
			elsif Bin = "00001101" then
			  x := "000000010011";
			elsif Bin = "1110" then
			  x := "000000010100";
			elsif Bin = "00001111" then
			  x := "000000010101";
			elsif Bin = "00010000" then
			  x := "000000010110";
			elsif Bin = "10001" then
			  x := "000000010111";
			elsif Bin = "00010010" then
			  x := "000000011000";
			elsif Bin = "00010011" then
			  x := "000000011001";
			elsif Bin = "00010100" then
			  x := "000000100000";
			elsif Bin = "00010101" then
			  x := "000000100001";
			elsif Bin = "00010110" then
			  x := "000000100010";
			elsif Bin = "10111" then
			  x := "000000100011";
			elsif Bin = "00011000" then
			  x := "000000100100";
			elsif Bin = "00011001" then
			  x := "000000100101";
			elsif Bin = "00011010" then
			  x := "000000100110";
			elsif Bin = "00011011" then
			  x := "000000100111";
			elsif Bin = "00011100" then
			  x := "000000101000";
			elsif Bin = "00011101" then
			  x := "000000101001";
			elsif Bin = "00011110" then
			  x := "000000110000";
			elsif Bin = "00011111" then
			  x := "000000110001";
			elsif Bin = "00100000" then
			  x := "000000110010";
			elsif Bin = "00100001" then
			  x := "000000110011";
			elsif Bin = "00100010" then
			  x := "000000110100";
			elsif Bin = "00100011" then
			  x := "000000110101";
			elsif Bin = "00100100" then
			  x := "000000110110";
			elsif Bin = "00100101" then
			  x := "000000110111";
			elsif Bin = "00100110" then
			  x := "000000111000";
			elsif Bin = "00100111" then
			  x := "000000111001";
			elsif Bin = "00101000" then
			  x := "000001000000";
			elsif Bin = "00101001" then
			  x := "000001000001";
			elsif Bin = "00101010" then
			  x := "000001000010";
			elsif Bin = "00101011" then
			  x := "000001000011";
			elsif Bin = "00101100" then
			  x := "000001000100";
			elsif Bin = "00101101" then
			  x := "000001000101";
			elsif Bin = "00101110" then
			  x := "000001000110";
			elsif Bin = "00101111" then
			  x := "000001000111";
			elsif Bin = "00110000" then
			  x := "000001001000";
			elsif Bin = "00110001" then
			  x := "000001001001";
			elsif Bin = "00110010" then
			  x := "000001010000";
			elsif Bin = "00110011" then
			  x := "000001010001";
			elsif Bin = "00110100" then
			  x := "000001010010";
			elsif Bin = "00110101" then
			  x := "000001010011";
			elsif Bin = "00110110" then
			  x := "000001010100";
			elsif Bin = "00110111" then
			  x := "000001010101";
			elsif Bin = "00111000" then
			  x := "000001010110";
			elsif Bin = "00111001" then
			  x := "000001010111";
			elsif Bin = "00111010" then
			  x := "000001011000";
			elsif Bin = "00111011" then
			  x := "000001011001";
			elsif Bin = "00111100" then
			  x := "000001100000";
			elsif Bin = "00111101" then
			  x := "000001100001";
			elsif Bin = "00111110" then
			  x := "000001100010";
			elsif Bin = "00111111" then
			  x := "000001100011";
			elsif Bin = "01000000" then
			  x := "000001100100";
			elsif Bin = "1000001" then
			  x := "000001100101";
			elsif Bin = "01000010" then
			  x := "000001100110";
			elsif Bin = "01000011" then
			  x := "000001100111";
			elsif Bin = "01000100" then
			  x := "000001101000";
			elsif Bin = "01000101" then
			  x := "000001101001";
			elsif Bin = "01000110" then
			  x := "000001110000";
			elsif Bin = "01000111" then
			  x := "000001110001";
			elsif Bin = "01001000" then
			  x := "000001110010";
			elsif Bin = "01001001" then
			  x := "000001110011";
			elsif Bin = "01001010" then
			  x := "000001110100";
			elsif Bin = "01001011" then
			  x := "000001110101";
			elsif Bin = "01001100" then
			  x := "000001110110";
			elsif Bin = "01001101" then
			  x := "000001110111";
			elsif Bin = "01001110" then
			  x := "000001111000";
			elsif Bin = "01001111" then
			  x := "000001111001";
			elsif Bin = "01010000" then
			  x := "000010000000";
			elsif Bin = "01010001" then
			  x := "000010000001";
			elsif Bin = "01010010" then
			  x := "000010000010";
			elsif Bin = "01010011" then
			  x := "000010000011";
			elsif Bin = "01010100" then
			  x := "000010000100";
			elsif Bin = "01010101" then
			  x := "000010000101";
			elsif Bin = "01010110" then
			  x := "000010000110";
			elsif Bin = "01010111" then
			  x := "000010000111";
			elsif Bin = "01011000" then
			  x := "000010001000";
			elsif Bin = "01011001" then
			  x := "000010001001";
			elsif Bin = "01011010" then
			  x := "000010010000";
			elsif Bin = "01011011" then
			  x := "000010010001";
			elsif Bin = "01011100" then
			  x := "000010010010";
			elsif Bin = "01011101" then
			  x := "000010010011";
			elsif Bin = "01011110" then
			  x := "000010010100";
			elsif Bin = "01011111" then
			  x := "000010010101";
			elsif Bin = "01100000" then
			  x := "000010010110";
			elsif Bin = "01100001" then
			  x := "000010010111";
			elsif Bin = "1100010" then
			  x := "000010011000";
			elsif Bin = "01100011" then
			  x := "000010011001";
			elsif Bin = "01100100" then
			  x := "000100000000";
			elsif Bin = "01100101" then
			  x := "000100000001";
			elsif Bin = "01100110" then
			  x := "000100000010";
			elsif Bin = "01100111" then
			  x := "000100000011";
			elsif Bin = "01101000" then
			  x := "000100000100";
			elsif Bin = "01101001" then
			  x := "000100000101";
			elsif Bin = "01101010" then
			  x := "000100000110";
			elsif Bin = "01101011" then
			  x := "000100000111";
			elsif Bin = "01101100" then
			  x := "000100001000";
			elsif Bin = "01101101" then
			  x := "000100001001";
			elsif Bin = "01101110" then
			  x := "000100010000";
			elsif Bin = "01101111" then
			  x := "000100010001";
			elsif Bin = "01110000" then
			  x := "000100010010";
			elsif Bin = "01110001" then
			  x := "000100010011";
			elsif Bin = "01110010" then
			  x := "000100010100";
			elsif Bin = "1110011" then
			  x := "000100010101";
			elsif Bin = "01110100" then
			  x := "000100010110";
			elsif Bin = "01110101" then
			  x := "000100010111";
			elsif Bin = "01110110" then
			  x := "000100011000";
			elsif Bin = "01110111" then
			  x := "000100011001";
			elsif Bin = "01111000" then
			  x := "000100100000";
			elsif Bin = "01111001" then
			  x := "000100100001";
			elsif Bin = "01111010" then
			  x := "000100100010";
			elsif Bin = "01111011" then
			  x := "000100100011";
			elsif Bin = "01111100" then
			  x := "000100100100";
			elsif Bin = "01111101" then
			  x := "000100100101";
			elsif Bin = "01111110" then
			  x := "000100100110";
			elsif Bin = "01111111" then
			  x := "000100100111";
			elsif Bin = "10000000" then
			  x := "000100101000";
			elsif Bin = "10000001" then
			  x := "000100101001";
			elsif Bin = "10000010" then
			  x := "000100110000";
			elsif Bin = "10000011" then
			  x := "000100110001";
			elsif Bin = "10000100" then
			  x := "000100110010";
			elsif Bin = "10000101" then
			  x := "000100110011";
			elsif Bin = "10000110" then
			  x := "000100110100";
			elsif Bin = "10000111" then
			  x := "000100110101";
			elsif Bin = "10001000" then
			  x := "000100110110";
			elsif Bin = "10001001" then
			  x := "000100110111";
			elsif Bin = "10001010" then
			  x := "000100111000";
			elsif Bin = "10001011" then
			  x := "000100111001";
			elsif Bin = "10001100" then
			  x := "000101000000";
			elsif Bin = "10001101" then
			  x := "000101000001";
			elsif Bin = "10001110" then
			  x := "000101000010";
			elsif Bin = "10001111" then
			  x := "000101000011";
			elsif Bin = "10010000" then
			  x := "000101000100";
			elsif Bin = "10010001" then
			  x := "000101000101";
			elsif Bin = "10010010" then
			  x := "000101000110";
			elsif Bin = "10010011" then
			  x := "000101000111";
			elsif Bin = "10010100" then
			  x := "000101001000";
			elsif Bin = "10010101" then
			  x := "000101001001";
			elsif Bin = "10010110" then
			  x := "000101010000";
			elsif Bin = "10010111" then
			  x := "000101010001";
			elsif Bin = "10011000" then
			  x := "000101010010";
			elsif Bin = "10011001" then
			  x := "000101010011";
			elsif Bin = "10011010" then
			  x := "000101010100";
			elsif Bin = "10011011" then
			  x := "000101010101";
			elsif Bin = "10011100" then
			  x := "000101010110";
			elsif Bin = "10011101" then
			  x := "000101010111";
			elsif Bin = "10011110" then
			  x := "000101011000";
			elsif Bin = "10011111" then
			  x := "000101011001";
			elsif Bin = "10100000" then
			  x := "000101100000";
			elsif Bin = "10100001" then
			  x := "000101100001";
			elsif Bin = "10100010" then
			  x := "000101100010";
			elsif Bin = "10100011" then
			  x := "000101100011";
			elsif Bin = "10100100" then
			  x := "000101100100";
			elsif Bin = "10100101" then
			  x := "000101100101";
			elsif Bin = "10100110" then
			  x := "000101100110";
			elsif Bin = "10100111" then
			  x := "000101100111";
			elsif Bin = "10101000" then
			  x := "000101101000";
			elsif Bin = "10101001" then
			  x := "000101101001";
			elsif Bin = "10101010" then
			  x := "000101110000";
			elsif Bin = "10101011" then
			  x := "000101110001";
			elsif Bin = "10101100" then
			  x := "000101110010";
			elsif Bin = "10101101" then
			  x := "000101110011";
			elsif Bin = "10101110" then
			  x := "000101110100";
			elsif Bin = "10101111" then
			  x := "000101110101";
			elsif Bin = "10110000" then
			  x := "000101110110";
			elsif Bin = "10110001" then
			  x := "000101110111";
			elsif Bin = "10110010" then
			  x := "000101111000";
			elsif Bin = "10110011" then
			  x := "000101111001";
			elsif Bin = "10110100" then
			  x := "000110000000";
			elsif Bin = "10110101" then
			  x := "000110000001";
			elsif Bin = "10110110" then
			  x := "000110000010";
			elsif Bin = "10110111" then
			  x := "000110000011";
			elsif Bin = "10111000" then
			  x := "000110000100";
			elsif Bin = "10111001" then
			  x := "000110000101";
			elsif Bin = "10111010" then
			  x := "000110000110";
			elsif Bin = "10111011" then
			  x := "000110000111";
			elsif Bin = "10111100" then
			  x := "000110001000";
			elsif Bin = "10111101" then
			  x := "000110001001";
			elsif Bin = "10111110" then
			  x := "000110010000";
			elsif Bin = "10111111" then
			  x := "000110010001";
			elsif Bin = "11000000" then
			  x := "000110010010";
			elsif Bin = "11000001" then
			  x := "000110010011";
			elsif Bin = "11000010" then
			  x := "000110010100";
			elsif Bin = "11000011" then
			  x := "000110010101";
			elsif Bin = "11000100" then
			  x := "000110010110";
			elsif Bin = "11000101" then
			  x := "000110010111";
			elsif Bin = "11000110" then
			  x := "000110011000";
			elsif Bin = "11000111" then
			  x := "000110011001";
			elsif Bin = "11001000" then
			  x := "001000000000";
			elsif Bin = "11001001" then
			  x := "001000000001";
			elsif Bin = "11001010" then
			  x := "001000000010";
			elsif Bin = "11001011" then
			  x := "001000000011";
			elsif Bin = "11001100" then
			  x := "001000000100";
			elsif Bin = "11001101" then
			  x := "001000000101";
			elsif Bin = "11001110" then
			  x := "001000000110";
			elsif Bin = "11001111" then
			  x := "001000000111";
			elsif Bin = "11010000" then
			  x := "001000001000";
			elsif Bin = "11010001" then
			  x := "001000001001";
			elsif Bin = "11010010" then
			  x := "001000010000";
			elsif Bin = "11010011" then
			  x := "001000010001";
			elsif Bin = "11010100" then
			  x := "001000010010";
			elsif Bin = "11010101" then
			  x := "001000010011";
			elsif Bin = "11010110" then
			  x := "001000010100";
			elsif Bin = "11010111" then
			  x := "001000010101";
			elsif Bin = "11011000" then
			  x := "001000010110";
			elsif Bin = "11011001" then
			  x := "001000010111";
			elsif Bin = "11011010" then
			  x := "001000011000";
			elsif Bin = "11011011" then
			  x := "001000011001";
			elsif Bin = "11011100" then
			  x := "001000100000";
			elsif Bin = "11011101" then
			  x := "001000100001";
			elsif Bin = "11011110" then
			  x := "001000100010";
			elsif Bin = "11011111" then
			  x := "001000100011";
			elsif Bin = "11100000" then
			  x := "001000100100";
			elsif Bin = "11100001" then
			  x := "001000100101";
			elsif Bin = "11100010" then
			  x := "001000100110";
			elsif Bin = "11100011" then
			  x := "001000100111";
			elsif Bin = "11100100" then
			  x := "001000101000";
			elsif Bin = "11100101" then
			  x := "001000101001";
			elsif Bin = "11100110" then
			  x := "001000110000";
			elsif Bin = "11100111" then
			  x := "001000110001";
			elsif Bin = "11101000" then
			  x := "001000110010";
			elsif Bin = "11101001" then
			  x := "001000110011";
			elsif Bin = "11101010" then
			  x := "001000110100";
			elsif Bin = "11101011" then
			  x := "001000110101";
			elsif Bin = "11101100" then
			  x := "001000110110";
			elsif Bin = "11101101" then
			  x := "001000110111";
			elsif Bin = "11101110" then
			  x := "001000111000";
			elsif Bin = "11101111" then
			  x := "001000111001";
			elsif Bin = "11110000" then
			  x := "001001000000";
			elsif Bin = "11110001" then
			  x := "001001000001";
			elsif Bin = "11110010" then
			  x := "001001000010";
			elsif Bin = "11110011" then
			  x := "001001000011";
			elsif Bin = "11110100" then
			  x := "001001000100";
			elsif Bin = "11110101" then
			  x := "001001000101";
			elsif Bin = "11110110" then
			  x := "001001000110";
			elsif Bin = "11110111" then
			  x := "001001000111";
			elsif Bin = "11111000" then
			  x := "001001001000";
			elsif Bin = "11111001" then
			  x := "001001001001";
			elsif Bin = "11111010" then
			  x := "001001010000";
			elsif Bin = "11111011" then
			  x := "001001010001";
			elsif Bin = "11111100" then
			  x := "001001010010";
			elsif Bin = "11111101" then
			  x := "001001010011";
			elsif Bin = "11111110" then
			  x := "001001010100";
			elsif Bin = "11111111" then 
			  x := "001001010101";
			end if;
        Cen <= x(11 downto 8);
        Dec <= x(7 downto 4);
        Uni <= x(3 downto 0);
    end process;
    
end Behavioral;