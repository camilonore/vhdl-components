library verilog;
use verilog.vl_types.all;
entity t_flipflop_vlg_vec_tst is
end t_flipflop_vlg_vec_tst;
