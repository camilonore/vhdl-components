library verilog;
use verilog.vl_types.all;
entity divisor_2_vlg_sample_tst is
    port(
        Clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end divisor_2_vlg_sample_tst;
